module tx_counter (input clk,
                   input reset,
                   input count_enable,
                   output reg count_out);

    reg [3:0] count;

    always @(posedge clk) begin
        count_out <= 0;
        if (!reset) begin
            count <= 0;
        end
        else if (count) begin
            if (count == 9) begin
                count <= 0;
                count_out <= 1;
            end
            else begin
                count <= count + 1;
            end
        end
    end
endmodule